amp application

*-----------------------------------------------------------------------------

V1 in 0 0.0 ac 1.0 SIN(1.65 10 1kHz)
r1 in vout 1k
*d1 n 0 d1n5913brl
*d2 n vout d1n5913brl
*d1 0 n CMDZ5226B
*d2 vout n CMDZ5226B

d1 0 vout Dbreak

.model Dbreak d Is=1e-14 Cjo=1e-11 Rs=0.1 BV=3.3v IBV=2mA

*-----------------------------------------------------------------------------
*SRC=CMDZ5226B;CMDZ5226B;Diodes;Zener <=10V; 3.30V  0.250W   CENTRAL -
*SYM=HZEN
.SUBCKT CMDZ5226B  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 0.716
.MODEL DF D ( IS=31.2p RS=2.56 N=1.10
+ CJO=270p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=6.24f RS=17.3 N=3.00 )
.ENDS
*-----------------------------------------------------------------------------
.SUBCKT d1n5913brl 2 1
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*    Modeling services provided by   *
* Interface Technologies www.i-t.com *
**************************************
* Model generated on Jun 22, 2004
* MODEL FORMAT: SPICE3
*     anode cathode
*node: 2      1
*    Forward Section
D1 2 1 MD1
.MODEL MD1 D IS=1.33275e-21 N=1 XTI=1 RS=0.1
+ CJO=1e-11 TT=1e-08
*    Leakage Current
R 1 2 10000 MDR	
.MODEL MDR R TC1=0 TC2=0
*    Breakdown
RZ 2 3 8.29777
IZG 4 3 0.5448
R4 4 3 500
D3 3 4 MD3
.MODEL MD3 D IS=2.5e-12 N=4.68677 XTI=0 EG=0.1
D2 5 4 MD2
.MODEL MD2 D IS=2.5e-12 N=6.25163 XTI=0 EG=0.1
EV1 1 5 6 0 1
IBV 0 6 0.001
RBV 6 0 1526.95 MDRBV
.MODEL MDRBV R TC1=-6.06e-08
*-- SPICE3 DIODE MODEL DEFAULT PARAMETER
*  VALUES ARE ASSUMED
*IS=1E-14 RS=0 N=1 TT=0 CJO=0
*VJ=1 M=0.5 EG=1.11 XTI=3 FC=0.5
*KF=0 AF=1 BV=inf IBV=1e-3 TNOM=27
.ENDS d1n5913brl
---------------------------------------------------------------

.control
  set hcopydevtype=postscript

* color0 is background color
* color1 is the grid and text color
* colors 2-15 are for the vectors if you want to specify them
* uncomment next three lines to plot colors on white background
  set hcopypscolor=true
  set color0=rgb:f/f/f
  set color1=rgb:0/0/0

* to print the results directly to a printer uncomment the following line
* set hcopydev=kec3112

* run DC operating point simulation first
  op

*run transient simulation for 40ns with timesteps of 100ps
  tran 1e-5 2e-3

*plot nodes tline_input and tline_output every 1ns for 45ns
  plot in vout

*plot to .ps file nodes tline_input and tline_output every 1ns for 45ns
 * hardcopy tline_plot.ps V(tline_input) V(tline_output) xl 0.1ns 40ns

.endc

.end
