amp application

*-----------------------------------------------------------------------------

V1 vin 0  0.0 ac 1.0 SIN(2.5 2.5 1Hz)
*V1 vin 0 dc 0.5
V2 v5v 0 dc 5
v3 v3v 0 dc 3.3
v4 vpwm 0 dc 1

*xor in rfg vcc 0 aout uA741
*xorb vrefi about vcc 0 about uA741
xor anin aiin v5v 0 aout LMC6032/NS
xorb aout bout v5v 0 bout LMC6032/NS

r1 vin anin 10k
r2 anin 0 36.5k
c1 vin 0 470pf
c2 anin 0 10uf
r3 aiin aout 10k
r4 aiin v5v 82.5k
r5 aiin 0 665k
r6 aiin m1 33.2k
r7 m1 vpwm 33.2k
c3 m1 0 1uf
r8 bout 0 1k
r9 bout n1 24k
r10 n1 n2 4k
r11 n2 n3 2k
r12 n3 n4 1k
r13 n4 0 2k
r14 n4 v3v 2k

*ddd1 0 vout Dbreak

*.model Dbreak d Is=1e-14 Cjo=1e-11 Rs=0.1 BV=3.3v IBV=2mA

*d1 0 vout d1n5913brl
*d1 0 vout CMDZ5226B



*-----------------------------------------------------------------------------
*SRC=CMDZ5226B;CMDZ5226B;Diodes;Zener <=10V; 3.30V  0.250W   CENTRAL -
*SYM=HZEN
.SUBCKT CMDZ5226B  1 2
*Terminals         A C
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 0.716
.MODEL DF D ( IS=31.2p RS=2.56 N=1.10
+ CJO=270p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=6.24f RS=17.3 N=3.00 )
.ENDS
*-----------------------------------------------------------------------------
.SUBCKT d1n5913brl 2 1
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*    Modeling services provided by   *
* Interface Technologies www.i-t.com *
**************************************
* Model generated on Jun 22, 2004
* MODEL FORMAT: SPICE3
*     anode cathode
*node: 2      1
*    Forward Section
D1 2 1 MD1
.MODEL MD1 D IS=1.33275e-21 N=1 XTI=1 RS=0.1
+ CJO=1e-11 TT=1e-08
*    Leakage Current
R 1 2 10000 MDR	
.MODEL MDR R TC1=0 TC2=0
*    Breakdown
RZ 2 3 8.29777
IZG 4 3 0.5448
R4 4 3 500
D3 3 4 MD3
.MODEL MD3 D IS=2.5e-12 N=4.68677 XTI=0 EG=0.1
D2 5 4 MD2
.MODEL MD2 D IS=2.5e-12 N=6.25163 XTI=0 EG=0.1
EV1 1 5 6 0 1
IBV 0 6 0.001
RBV 6 0 1526.95 MDRBV 
.MODEL MDRBV R TC1=-6.06e-08
*-- SPICE3 DIODE MODEL DEFAULT PARAMETER
*  VALUES ARE ASSUMED
*IS=1E-14 RS=0 N=1 TT=0 CJO=0
*VJ=1 M=0.5 EG=1.11 XTI=3 FC=0.5
*KF=0 AF=1 BV=inf IBV=1e-3 TNOM=27
.ENDS d1n5913brl


*-----------------------------------------------------------------------------
* To use a subcircuit, the name must begin with 'X'.  For example:
* X1 1 2 3 4 5 uA741
*
* connections:   non-inverting input
*                |  inverting input
*                |  |  positive power supply
*                |  |  |  negative power supply
*                |  |  |  |  output
*                |  |  |  |  |
.subckt uA741    1  2  3  4  5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*-----------------------------------------------------------------------------
* LMC6032 CMOS Dual Operational Amplifier
* ////////////////////////////////////////
*
* Connections:      Non-inverting input
*                   |   Inverting input
*                   |   |   Positive power supply
*                   |   |   |   Negative power supply
*                   |   |   |   |   Output
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LMC6032/NS  1   2  99  50  28
* CAUTION:  SET .OPTIONS GMIN=1E-16 TO CORRECTLY MODEL INPUT BIAS CURRENT.
*
* Features:
* Operates from single supply
* Rail-to-rail output swing
* Low offset voltage (max) =             9mV
* Ultra low input current =              2fA
* Slew rate =                        1.1V/uS
* Gain-bandwidth product =           1.4 MHz 
* Low supply current =                 375uA/Amplifier
*
* NOTE: - Model is for single device only and simulated
*         supply current is 1/2 of total device current.
*       - Noise is not modeled.
*       - Asymmetrical gain is not modeled.
*
CI1 1  50 2P
CI2 2  50 2P
* 1.4 Hz pole capacitor
C3  98 9  11.35N
* 2.95 MHz pole capacitor
C4  6  5  4.93P
* Drain-substrate capacitor
C6  50 4  10P
* 35 MHz pole capacitor
C7  98 11 4.54F
DP1 1  99 DA
DP2 50 1  DX
DP3 2  99 DB
DP4 50 2  DX
D1  9  8  DX
D2  10 9  DX
D3  15 20 DX
D4  21 15 DX
D5  26 24 DX
D6  25 27 DX
D7  22 99 DX
D8  50 22 DX
D9  0  14 DX
D10 12 0  DX
EH  97 98 99    49 1.0
EN  0  96 0     50 1.0
* Input offset voltage -|
EOS 7  1  POLY(1) 16 49 9M 1
EP  97 0  99    0  1.0
E1  97 19 99    15 1.0
* Sourcing load +Vs current
F1  99 0  VA2   1
* Sinking load -Vs current
F2  0  50 VA3   1
F3  13 0  VA1   1
G1  98 9  5     6  0.1
G2  98 11 9     49 1U
G3  98 15 11    49 1U
* DC CMRR
G4  98 16 POLY(2) 1 49 2 49 0 3.54E-8 3.54E-8
I1  99 4  48.19U
I2  99 50 308.1U
* Load dependent pole
L1  22 28 40.4U
* CMR lead
L2  16 17 7.95M
M1  5  2  4     99 MX
M2  6  7  4     99 MX
R3  5  50 5.47K
R4  6  50 5.47K
R5  98 9  1E7
R8  99 49 133.3K
R9  49 50 133.3K
R12 98 11 1E6
R13 98 17 1K
* -Rout
R16 23 24 75
* +Rout
R17 23 25 70
* +Isc slope control
R18 20 29 144.6K
* -Isc slope control
R19 21 30 185K
R21 98 15 1E6
R22 22 28 900
VA1 19 23 0V
VA2 14 13 0V
VA3 13 12 0V
V2  97 8  0.721V
V3  10 96 0.721V
V4  29 22 0.63V
V5  22 30 0.63V
V6  26 22 0.63V
V7  22 27 0.63V
.MODEL  DA D    (IS=1.3E-14)
.MODEL  DB D    (IS=1.2E-14)
.MODEL  DX D    (IS=1.0E-14)
.MODEL  MX PMOS (VTO=-2.45 KP=7.0547E-4)
.ENDS

*-----------------------------------------------------------------------------

.control
  set hcopydevtype=postscript

* color0 is background color
* color1 is the grid and text color
* colors 2-15 are for the vectors if you want to specify them
* uncomment next three lines to plot colors on white background
  set hcopypscolor=true
  set color0=rgb:f/f/f
  set color1=rgb:0/0/0

* to print the results directly to a printer uncomment the following line
* set hcopydev=kec3112

* run DC operating point simulation first
  op

*run transient simulation for 40ns with timesteps of 100ps
  tran 1e-2 2e-0

*plot nodes tline_input and tline_output every 1ns for 45ns
  plot vin bout

*plot to .ps file nodes tline_input and tline_output every 1ns for 45ns
 * hardcopy tline_plot.ps V(tline_input) V(tline_output) xl 0.1ns 40ns

.endc

.end
